module ROB (
input clk,rst,write,
input [4:0] dest_reg, val_idx,
input [31:0] value,
output [4:0] tag,
output reg [4:0] commit_addr,
output reg [31:0] commit_val,
output reg full
);

reg [4:0] dest_regs [31:0];
reg [31:0] values [31:0];
reg [31:0] ready;
reg [4:0] issue_p,commit_p;


assign tag = issue_p;

always @(posedge clk, negedge rst) begin
	integer i;
	full = issue_p[3:0] + 1 == commit_p;
	if (~rst) begin
		ready = 0;
		issue_p=0;
		commit_p=0;
		for(i=0; i<32; i = i + 1) begin
			dest_regs[i] = 0;
			values[i] = 0;
		end
	end
	else begin
		if(~full) begin 
			dest_regs[issue_p] = dest_reg;
			ready[issue_p] = 0;
			issue_p = issue_p + 5'b1;
		end
		if (write) begin
			values[val_idx] = value;
			ready[val_idx] = 1;
		end
		if (ready[commit_p] == 1) begin
			commit_addr = dest_regs[commit_p];
			commit_val = values [commit_p];
			commit_p = commit_p +5'b1;		
		end
		
		
	end
	

end




endmodule