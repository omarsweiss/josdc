module retardmemory(clk,address,instruction);
	input clk;
	input [9:0] address;
	output reg [31:0] instruction;
	reg [31:0] data [1023:0];
	initial 
		begin
			data[0] = 32'b00100000000010000000000000001010;
data[1] = 32'b00100000000010010000000000010100;
data[2] = 32'b00000001000010010101000000100000;
data[3] = 32'b00000001001010000101100000100010;
data[4] = 32'b00000001000010010110000000100100;
data[5] = 32'b00000001000010010110100000100101;
data[6] = 32'b00000001000010010111000000100111;
data[7] = 32'b00000001000010010111100000100110;
data[8] = 32'b00100001000110000000000000001010;
data[9] = 32'b00110101001110010000000000000101;
data[10] = 32'b00111001001100000000000000000011;
data[11] = 32'b00000001000010011000100000101010;
data[12] = 32'b00000001000000001001000010000000;
data[13] = 32'b00000001001000001001100001000010;
data[14] = 32'b10101100000010100000000000000100;
data[15] = 32'b10001100000010110000000000000100;
data[16] = 32'b00010001001010000000000000000001;
data[17] = 32'b00010101001010000000000000000010;
data[18] = 32'b00100000000001000000000000000001;
data[19] = 32'b00001000000000000000000000011001;
data[20] = 32'b00100000000001000000000000000010;
data[21] = 32'b00001100000000000000000000010111;
data[22] = 32'b00001000000000000000000000011001;
data[23] = 32'b00100000000000100000000000000100;
data[24] = 32'b00000011111000000000000000000000;
data[25] = 32'b00100000000010000000000000000000;
end
	always @ (posedge clk)
		begin
			instruction = data[address];
		end


endmodule			